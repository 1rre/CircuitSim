*Netlist
V1 N001 0 SINE(0.75 1 1k)
R1 N002 N001 5k
R3 N003 0 16k
L1 N002 N003 100p
.tran 0 10m
.end
