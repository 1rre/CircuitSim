*Netlist
V1 N001 0 EXP(-2 5 450u 1.5m 6m 260u)
R1 N002 N001 5k
C3 N003 N002 160p
R1 N003 0 9.4k
.tran 0 10m
.end
