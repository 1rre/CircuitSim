*Netlist
V1 N001 0 SINE(50m 1.67 245 4.6m 100 795.4m 8)
R1 N003 N002 5k
R3 N004 0 16k
R2 N003 N004 3.2k
R4 N004 N003 0.032Meg
V3 N001 N002 PULSE(300m -400m 2m 1.9m 3.1m 500u 7.5m 5)
R5 N003 0 1Meg
R6 N004 N005 100k
V2 N003 N005 SFFM(0.0 1.6 4k 1.5 1.50k)
R7 N005 0 30k
.tran 0 50m
.end
