*Netlist
R1 N001 N002 5k
L3 N002 N003 160n
R1 N003 0 9.4k
V1 N001 0 EXP(2 5 450u 1.5m 6m 260u)
.tran 0 10m
.end
